IL is 10ma, find IV (Rs=0 , Rsh=5000)



*two diode equivalent of a solar cell
.subckt tdeq_solarcell IN OUT
rs IN 1 0
rsh 1 OUT 5000
d2 1 OUT diode2
.model diode2 d (is=(2e-6) n=2)
d1 1 OUT diode
.model diode d (is=(1e-13) n=1)
ic OUT 1 0.01
.ends

X1 2 0 tdeq_solarcell
vsource 1 0 dc 2
ra 1 2 100


.dc vsource -2 2 0.1

.control
run
plot  {(v(2)-v(1))*0.01} vs {v(2)}
.endc
.end
