RC Circuits


r1 2 3 1000
c1 3 0 1u
vin 2 0 pwl (0 -5v 0.005 -5v 0.0051 5v 0.01 5v 0.015) r=0

.control
*tran 0.01 0.35
*plot v(2)
*plot v(3)
*plot v(2) vs v(3)
*plot v(2) and v(3)
plot v(2) v(3)
plot v(2)
.endc
.end