RC Circuit with square wave with offset duty cycle 10% f=100Hz tran 0.0001m 30m


r1 2 3 1000
c1 3 0 1u
.param f = 100
.param width = {0.05/f}
.param period = {1/f}

vin 1 0 pulse(-5 5 0ns 0ns 0ns width period)
voffset 2 1 dc 5v
.control
run
tran 0.0001m 30m
plot v(2)v(3)
.endc
.end
