RC Q3 freequency response


r1 2 3 1000
c1 3 0 1u
vin 2 0 dc 0 ac 1

.ac dec 10 50 50000

.control 
run
plot vdb(3) xlog
plot {57.29*vp(3)} xlog 
plot vdb(3) {57.29*vp(3)} xlog 

.endc
.end
