I-V Characteristics of CD4007
.include cd4007.txt
vgg 1 0 dc 3.5v
rg 1 2 680
m1 3 2 0 0 NMOS4007
rd 3 4 100
vid 5 4 dc 0v
vdd 5 0 dc 0v
*Fixing Vgg, and varying Vdd from 0 to 5 in each case
.dc vdd 0 5 0.01 vgg 1 5 1
.control
run
plot vid#branch
.endc
.end
