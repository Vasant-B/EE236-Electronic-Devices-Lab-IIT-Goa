IL is 10ma, find IV (Rs=0 , Rsh=100)



*two diode equivalent of a solar cell
.subckt tdeq_solarcell IN OUT rs=0 rsh=100 ic=1
rs IN 1 {rs}
rsh 1 OUT {rsh}
d2 1 OUT diode2
.model diode2 d (is=(2e-6) n=2)
d1 1 OUT diode
.model diode d (is=(1e-13) n=1)
ic OUT 1 {ic}
.ends

X1 2 0 tdeq_solarcell rs=0 rsh=100 ic=0.01
vsource 1 0 dc 2
ra 1 2 100


.dc vsource -2 2 0.1
.control
run
plot  {(v(2)-v(1))*0.01} vs v(2)
.endc
.end

