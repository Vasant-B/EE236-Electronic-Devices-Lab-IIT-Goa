RC Circuits (without Log)


r1 2 3 1000
c1 3 0 1u
vin 2 0 dc 0 ac 1
.ac lin 100 50 50000
.control 
run
*tran 0.02m 0.35
*plot v(2)
plot v(3)
*plot v(2) vs v(3)
*plot v(2) and v(3)
*plot v(2) v(3)
plot vdb(3) xlog
plot {57.29*vp(3)} 
.endc
.end



*depratim sirs ppt
*RC Circuit Frequency Response 
*r1 1 2 1k 
*c1 2 0 1u 
*Specifying an AC source with zero dc 
*vin 1 0 dc 0 ac 1 
*AC analysis for 1 Hz to 1MHz, 10 points per decade 
*.ac dec 10 1 1Meg 
*.control 
*run 
*Magnitude dB plot for v(2) on log scale 
*plot vdb(2) xlog 
*Phase degrees plot for v(2) on log scale 
*plot {57.29*vp(2)} xlog 
*.endc 
*.end