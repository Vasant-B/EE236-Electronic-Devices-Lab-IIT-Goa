q6

.model bc547b NPN BF=500 NE=1.3 ISE=9.72F IKF=80M IS=20F 
+ VAF=50 ikr=12m BR=10 NC=2 VAR=10 RB=280 RE=1 RC=40 
+ VJE=.48 tr=.3u tf=.5n cje=12p vje=.48 mje=.5 cjc=6p 
+ vjc=.7 mjc=.33 isc=47p kf=2f

q1 3 7 2 bc547b
re 1 0 2000
rc 5 4 3000
r1 5 6 27000
r2 6 0 10000
vammeter_e 2 1 0
vammeter_c 4 3 0
vammeter_b 6 7 0
vcc 5 0 10v
vin 8 0 dc 0 ac 1
*sin(0 10m 5k 0 0)
cb 8 6 10mf
ce 1 0 10mf
cc 3 9 10mf
rl 9 0 1k

*AC analysis for 1 Hz to 1MHz, 10 points per decade 
.ac dec 10 1 1Meg 
.control 
run 
*Magnitude dB plot for v(2) on log scale 
plot vdb(2) xlog 

*Phase degrees plot for v(2) on log scale 
plot {57.29*vp(2)} xlog 

*.tran 0.001m 2m
*.control
*run
*plot v(8) v(9)
*.endc
*.end