RC Q1 Vin=10Vpp 50Hz sine, r=1k, c=1u


r1 2 3 1000
c1 3 0 1u
vin 2 0 sin (0 5 50 0 0)

.control
tran 0.02m 0.35
plot v(2) v(3)
.endc
.end