CR Circuit with square wave  with offset


r1 3 0 1000
c1 2 3 1u
.param f = 100
.param width = {0.5/f}
.param period = {1/f}

vin 1 0 pulse(-5 5 0ns 0ns 0ns width period)
voffset 2 1 dc 5v
.control
run
tran 0.05m 100m
plot v(2)v(3)
.endc
.end
