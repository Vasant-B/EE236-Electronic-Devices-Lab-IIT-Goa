q1

.include BC547.txt

q1 1 2 3 bc547b
vce 1 3 5v
ic 1 4 1
vcc 0 4 10
vam1 3 0 0
r2 2 0 10k


.control
run
print v(2)
print vam#branch
.endc
.end