RC Circuit with square wave f(hz)=50,000 tran 0.001m 5m


r1 1 2 1000
c1 2 0 1u
.param f = 50000
.param width = {0.5/f}
.param period = {1/f}

vin 1 0 pulse(-5 5 0ns 0ns 0ns width period)

.control
run
tran 0.001m 5m
plot v(1)v(2)
.endc
.end
